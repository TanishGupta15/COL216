LIBRARY IEEE;
    USE IEEE.STD_LOGIC_1164.ALL;
    USE IEEE.STD_LOGIC_UNSIGNED.ALL;


--Only halt the program when special instruction HALT is received and not when instruction 0 is recieved.

ENTITY testbench IS 
-- empty
END ENTITY;

ARCHITECTURE BEV OF testbench IS


signal clk: std_logic;
signal input: std_logic_vector(7 downto 0);
signal status_bit: std_logic;
signal reset: std_logic;

-- DUT component
COMPONENT processor IS
    port (
    
    	clk: in std_logic;
		input: in std_logic_vector(7 downto 0);
		status_bit: in std_logic;
		reset: in std_logic;
    );
END COMPONENT;

BEGIN

  -- Connect DUT
  DUT: processor PORT MAP(
  clk => clk,
  input => input,
  status_bit => status_bit,
  reset => reset
  );

  PROCESS
  BEGIN
  	reset <= '0';
    status_bit <= '0';
    input <= X"00";
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
     wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
        wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
     wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
        wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
     wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
        wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
     wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
        wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
     wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
        wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
     wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
        wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
     wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
        wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
     wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
        wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
     wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
        wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
     wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
        wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
     wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
        wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
     wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
        wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
     wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
        wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
     wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
        wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
     wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
        wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
     wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
        wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
     wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
        wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
     wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
        wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
     wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
        wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
     wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
        wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
     wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
        wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
     wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
        wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
     wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
        wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
     wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
        wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
     wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
        wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
     wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
        wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
     wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
        wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
     wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
        wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
     wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
        wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
     wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
        wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
     wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
        wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    input <= X"24";
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    status_bit <= '1';
     wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
        wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
     wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
        wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
     wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
        wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
     wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    status_bit <= '0';
        wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
     wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
        wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
     wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
        wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
     wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
        wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
     wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
        wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
     wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
        wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
     wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
        wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1'; wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
        wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
     wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
        wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait for 1 ns;
    clk <= '0';
    wait for 1 ns;
    clk <= '1';
    wait;
  END PROCESS;

END BEV;
